library IEEE;
use IEEE.std_logic_1164.ALL;

entity flipflop is
   port(clk : in  std_logic;
        d   : in  std_logic;
        q   : out  std_logic);
end flipflop;



