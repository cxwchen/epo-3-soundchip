configuration adder_9x9_behavioral_cfg of adder_9x9 is
   for behavioral
   end for;
end adder_9x9_behavioral_cfg;
