library IEEE;
use IEEE.std_logic_1164.ALL;

entity var_shift is
   port(Sel_Out   : in  std_logic_vector(7 downto 0);
        vel       : in  std_logic_vector(6 downto 0);
        Shift_Out : out std_logic_vector(6 downto 0));
end var_shift;

