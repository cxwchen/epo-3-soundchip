configuration adder_7x7_behavioral_cfg of adder_7x7 is
   for behavioral
   end for;
end adder_7x7_behavioral_cfg;
