configuration adder6x5_behavioral_cfg of adder6x5 is
   for behavioral
   end for;
end adder6x5_behavioral_cfg;
