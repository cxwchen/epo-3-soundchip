library IEEE;
use IEEE.std_logic_1164.ALL;

entity channel_op_tb is
end channel_op_tb;

