configuration vel_shifter_behavioral_cfg of vel_shifter is
   for behavioral
   end for;
end vel_shifter_behavioral_cfg;
