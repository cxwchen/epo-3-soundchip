library IEEE;
use IEEE.std_logic_1164.ALL;

entity seq_mult_tb is
end seq_mult_tb;

