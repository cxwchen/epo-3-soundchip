library IEEE;
use IEEE.std_logic_1164.ALL;

entity midi_decoder_tb is
end midi_decoder_tb;

