library IEEE;
use IEEE.std_logic_1164.ALL;

entity inputbuffer is
   port(clk : in  std_logic;
        d   : in  std_logic;
        q   : out  std_logic);
end inputbuffer;


