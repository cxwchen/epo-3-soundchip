library IEEE;
use IEEE.std_logic_1164.ALL;

architecture behavioral of vel_shfiter is
begin



end behavioral;

