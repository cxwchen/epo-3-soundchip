library IEEE;
use IEEE.std_logic_1164.ALL;

entity pwm_math_tb is
end pwm_math_tb;

