configuration adder_6x6_behavioral_cfg of adder_6x6 is
   for behavioral
   end for;
end adder_6x6_behavioral_cfg;
