library library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity inputbuffer is
    port (

    );
end entity inputbuffer;

architecture structural of inputbuffer is
    
begin
    

    
end architecture structural;
