library library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity counter is
    port (
        
    );
end entity counter;

architecture structural of counter is
    
begin
    
    
    
end architecture structural;