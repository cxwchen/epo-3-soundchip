configuration input_sel_behavioral_cfg of input_sel is
   for behavioral
   end for;
end input_sel_behavioral_cfg;
