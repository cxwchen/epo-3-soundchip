configuration pwm_math_synthesised_cfg of pwm_math is
   for synthesised
      -- skipping oai211d0bwp7t because it is not a local entity
      -- skipping aoi221d0bwp7t because it is not a local entity
      -- skipping oai221d0bwp7t because it is not a local entity
      -- skipping oai22d0bwp7t because it is not a local entity
      -- skipping aoi31d0bwp7t because it is not a local entity
      -- skipping ao32d0bwp7t because it is not a local entity
      -- skipping aoi32d0bwp7t because it is not a local entity
      -- skipping moai22d0bwp7t because it is not a local entity
      -- skipping aoi222d0bwp7t because it is not a local entity
      -- skipping invd0bwp7t because it is not a local entity
      -- skipping inr3d0bwp7t because it is not a local entity
      -- skipping oai21d0bwp7t because it is not a local entity
      -- skipping aoi22d0bwp7t because it is not a local entity
      -- skipping cknd1bwp7t because it is not a local entity
      -- skipping ao21d0bwp7t because it is not a local entity
      -- skipping nd2d0bwp7t because it is not a local entity
      -- skipping nr2d0bwp7t because it is not a local entity
      -- skipping ao221d0bwp7t because it is not a local entity
      -- skipping nd3d0bwp7t because it is not a local entity
      -- skipping oai32d0bwp7t because it is not a local entity
      -- skipping ind3d0bwp7t because it is not a local entity
      -- skipping nr3d0bwp7t because it is not a local entity
      -- skipping maoi22d0bwp7t because it is not a local entity
      -- skipping invd1bwp7t because it is not a local entity
      -- skipping ind2d0bwp7t because it is not a local entity
      -- skipping ioa21d0bwp7t because it is not a local entity
      -- skipping inr2d0bwp7t because it is not a local entity
      -- skipping an2d1bwp7t because it is not a local entity
      -- skipping fa1d0bwp7t because it is not a local entity
      -- skipping maoi222d0bwp7t because it is not a local entity
      -- skipping ha1d0bwp7t because it is not a local entity
      -- skipping aoi21d0bwp7t because it is not a local entity
      -- skipping buffd4bwp7t because it is not a local entity
   end for;
end pwm_math_synthesised_cfg;
