configuration var_shift_behavioral_rounding_cfg of var_shift is
   for behavioral_rounding
   end for;
end var_shift_behavioral_rounding_cfg;
