library library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity register is
    port (
        
        );
end entity register;

architecture structural of register is
    
begin
    
    
    
end architecture structural;
