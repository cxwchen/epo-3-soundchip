library library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity fsm is
    port (
        
        );
end entity fsm;

architecture structural of fsm is
    
begin
    
    
    
end architecture structural;
