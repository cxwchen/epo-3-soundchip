configuration adder6x5_synthesised_cfg of adder6x5 is
   for synthesised
      -- skipping ckxor2d4bwp7t because it is not a local entity
      -- skipping nd2d4bwp7t because it is not a local entity
      -- skipping nd2d0bwp7t because it is not a local entity
      -- skipping ind3d0bwp7t because it is not a local entity
      -- skipping nr2d0bwp7t because it is not a local entity
      -- skipping ind2d0bwp7t because it is not a local entity
      -- skipping oai211d0bwp7t because it is not a local entity
      -- skipping inr2d0bwp7t because it is not a local entity
      -- skipping oai21d0bwp7t because it is not a local entity
      -- skipping ckan2d4bwp7t because it is not a local entity
      -- skipping or2d0bwp7t because it is not a local entity
      -- skipping cknd2d1bwp7t because it is not a local entity
      -- skipping inr2d1bwp7t because it is not a local entity
      -- skipping invd4bwp7t because it is not a local entity
      -- skipping invd1bwp7t because it is not a local entity
   end for;
end adder6x5_synthesised_cfg;
