configuration seq_mult_behavioral_cfg of seq_mult is
   for behavioral
   end for;
end seq_mult_behavioral_cfg;
