configuration mult_adder_behavioral_cfg of mult_adder is
   for behavioral
   end for;
end mult_adder_behavioral_cfg;
