library IEEE;
use IEEE.std_logic_1164.ALL;

entity partial_mult_tb is
end partial_mult_tb;

