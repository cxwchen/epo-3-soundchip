configuration adder5x4_behavioral_cfg of adder5x4 is
   for behavioral
   end for;
end adder5x4_behavioral_cfg;
