configuration channel_adder_behavioral_cfg of channel_adder is
   for behavioral
   end for;
end channel_adder_behavioral_cfg;
