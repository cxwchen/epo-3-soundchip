configuration adder_8x8_behavioral_cfg of adder_8x8 is
   for behavioral
   end for;
end adder_8x8_behavioral_cfg;
