library IEEE;
use IEEE.std_logic_1164.ALL;

entity input_sel_tb is
end input_sel_tb;

