configuration var_shift_behavioral_cfg of var_shift is
   for behavioral
   end for;
end var_shift_behavioral_cfg;
